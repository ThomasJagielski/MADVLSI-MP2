magic
tech sky130A
timestamp 1614454945
<< nwell >>
rect -70 640 255 1395
<< nmos >>
rect 0 420 15 520
rect 40 420 55 520
rect 105 420 120 520
rect 170 420 185 520
rect 0 -65 15 35
rect 40 -65 55 35
rect 105 -65 120 35
rect 170 -65 185 35
<< pmos >>
rect 0 1140 15 1240
rect 65 1140 80 1240
rect 130 1140 145 1240
rect 170 1140 185 1240
rect 0 660 15 760
rect 65 660 80 760
rect 130 660 145 760
rect 170 660 185 760
<< ndiff >>
rect -50 505 0 520
rect -50 435 -35 505
rect -15 435 0 505
rect -50 420 0 435
rect 15 420 40 520
rect 55 505 105 520
rect 55 435 70 505
rect 90 435 105 505
rect 55 420 105 435
rect 120 505 170 520
rect 120 435 135 505
rect 155 435 170 505
rect 120 420 170 435
rect 185 505 235 520
rect 185 435 200 505
rect 220 435 235 505
rect 185 420 235 435
rect -50 20 0 35
rect -50 -50 -35 20
rect -15 -50 0 20
rect -50 -65 0 -50
rect 15 -65 40 35
rect 55 20 105 35
rect 55 -50 70 20
rect 90 -50 105 20
rect 55 -65 105 -50
rect 120 20 170 35
rect 120 -50 135 20
rect 155 -50 170 20
rect 120 -65 170 -50
rect 185 20 235 35
rect 185 -50 200 20
rect 220 -50 235 20
rect 185 -65 235 -50
<< pdiff >>
rect -50 1225 0 1240
rect -50 1155 -35 1225
rect -15 1155 0 1225
rect -50 1140 0 1155
rect 15 1225 65 1240
rect 15 1155 30 1225
rect 50 1155 65 1225
rect 15 1140 65 1155
rect 80 1225 130 1240
rect 80 1155 95 1225
rect 115 1155 130 1225
rect 80 1140 130 1155
rect 145 1140 170 1240
rect 185 1225 235 1240
rect 185 1155 200 1225
rect 220 1155 235 1225
rect 185 1140 235 1155
rect -50 745 0 760
rect -50 675 -35 745
rect -15 675 0 745
rect -50 660 0 675
rect 15 745 65 760
rect 15 675 30 745
rect 50 675 65 745
rect 15 660 65 675
rect 80 745 130 760
rect 80 675 95 745
rect 115 675 130 745
rect 80 660 130 675
rect 145 660 170 760
rect 185 745 235 760
rect 185 675 200 745
rect 220 675 235 745
rect 185 660 235 675
<< ndiffc >>
rect -35 435 -15 505
rect 70 435 90 505
rect 135 435 155 505
rect 200 435 220 505
rect -35 -50 -15 20
rect 70 -50 90 20
rect 135 -50 155 20
rect 200 -50 220 20
<< pdiffc >>
rect -35 1155 -15 1225
rect 30 1155 50 1225
rect 95 1155 115 1225
rect 200 1155 220 1225
rect -35 675 -15 745
rect 30 675 50 745
rect 95 675 115 745
rect 200 675 220 745
<< psubdiff >>
rect 15 -110 65 -95
rect 15 -180 30 -110
rect 50 -180 65 -110
rect 15 -195 65 -180
rect 120 -110 170 -95
rect 120 -180 135 -110
rect 155 -180 170 -110
rect 120 -195 170 -180
<< nsubdiff >>
rect 15 1355 65 1370
rect 15 1285 30 1355
rect 50 1285 65 1355
rect 15 1270 65 1285
rect 120 1355 170 1370
rect 120 1285 135 1355
rect 155 1285 170 1355
rect 120 1270 170 1285
<< psubdiffcont >>
rect 30 -180 50 -110
rect 135 -180 155 -110
<< nsubdiffcont >>
rect 30 1285 50 1355
rect 135 1285 155 1355
<< poly >>
rect 0 1240 15 1255
rect 65 1240 80 1255
rect 130 1240 145 1255
rect 170 1240 185 1255
rect 0 955 15 1140
rect 65 1085 80 1140
rect 130 1130 145 1140
rect 40 1075 80 1085
rect 40 1055 50 1075
rect 70 1055 80 1075
rect 40 1045 80 1055
rect 105 1115 145 1130
rect 170 1130 185 1140
rect 170 1115 200 1130
rect 40 1010 80 1020
rect 40 990 50 1010
rect 70 990 80 1010
rect 40 980 80 990
rect 0 940 40 955
rect 25 790 40 940
rect 0 775 40 790
rect 0 760 15 775
rect 65 760 80 980
rect 105 785 120 1115
rect 185 915 200 1115
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 105 770 145 785
rect 130 760 145 770
rect 170 760 185 810
rect 0 520 15 660
rect 65 650 80 660
rect 130 650 145 660
rect 40 635 80 650
rect 105 635 145 650
rect 40 520 55 635
rect 105 520 120 635
rect 170 520 185 660
rect 0 235 15 420
rect 40 365 55 420
rect 40 355 80 365
rect 40 335 50 355
rect 70 335 80 355
rect 40 325 80 335
rect 40 290 80 300
rect 40 270 50 290
rect 70 270 80 290
rect 40 260 80 270
rect 0 220 40 235
rect 25 100 40 220
rect 0 85 40 100
rect 0 35 15 85
rect 65 60 80 260
rect 40 45 80 60
rect 40 35 55 45
rect 105 35 120 420
rect 170 195 185 420
rect 170 185 225 195
rect 170 165 195 185
rect 215 165 225 185
rect 170 155 225 165
rect 145 120 185 130
rect 145 100 155 120
rect 175 100 185 120
rect 145 90 185 100
rect 170 35 185 90
rect 0 -210 15 -65
rect 40 -80 55 -65
rect 105 -210 120 -65
rect 170 -80 185 -65
rect -25 -220 15 -210
rect -25 -240 -15 -220
rect 5 -240 15 -220
rect -25 -245 15 -240
rect 80 -220 120 -210
rect 80 -240 90 -220
rect 110 -240 120 -220
rect 80 -245 120 -240
<< polycont >>
rect 50 1055 70 1075
rect 50 990 70 1010
rect 195 885 215 905
rect 155 820 175 840
rect 50 335 70 355
rect 50 270 70 290
rect 195 165 215 185
rect 155 100 175 120
rect -15 -240 5 -220
rect 90 -240 110 -220
<< locali >>
rect 20 1355 60 1365
rect 20 1285 30 1355
rect 50 1285 60 1355
rect 20 1275 60 1285
rect 125 1355 165 1365
rect 125 1285 135 1355
rect 155 1285 165 1355
rect 125 1275 165 1285
rect -50 1225 -5 1235
rect -50 1155 -35 1225
rect -15 1155 -5 1225
rect -50 1145 -5 1155
rect 20 1225 60 1235
rect 20 1155 30 1225
rect 50 1155 60 1225
rect 20 1145 60 1155
rect 85 1225 125 1235
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 1145 125 1155
rect 190 1225 235 1235
rect 190 1155 200 1225
rect 220 1155 235 1225
rect 190 1145 235 1155
rect 40 1125 60 1145
rect 190 1125 210 1145
rect 40 1105 120 1125
rect 40 1075 80 1085
rect 40 1065 50 1075
rect 0 1055 50 1065
rect 70 1055 80 1075
rect 0 1045 80 1055
rect 0 960 20 1045
rect 100 1020 120 1105
rect 40 1010 120 1020
rect 40 990 50 1010
rect 70 1000 120 1010
rect 145 1105 210 1125
rect 70 990 80 1000
rect 40 980 80 990
rect 0 940 40 960
rect 20 755 40 940
rect 145 850 165 1105
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 205 755 225 875
rect -50 745 -5 755
rect -50 675 -35 745
rect -15 675 -5 745
rect -50 665 -5 675
rect 20 745 60 755
rect 20 675 30 745
rect 50 675 60 745
rect 20 665 60 675
rect 85 745 125 755
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect 190 745 235 755
rect 190 675 200 745
rect 220 675 235 745
rect 190 665 235 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect 40 515 60 665
rect 190 640 210 665
rect 145 620 210 640
rect 145 515 165 620
rect 40 505 100 515
rect 40 495 70 505
rect -50 425 -5 435
rect 60 435 70 495
rect 90 435 100 505
rect 60 425 100 435
rect 125 505 165 515
rect 125 435 135 505
rect 155 435 165 505
rect 125 425 165 435
rect 190 505 235 515
rect 190 435 200 505
rect 220 435 235 505
rect 190 425 235 435
rect 80 405 100 425
rect 80 385 120 405
rect 40 355 80 365
rect 40 345 50 355
rect 0 335 50 345
rect 70 335 80 355
rect 0 325 80 335
rect 0 240 20 325
rect 100 300 120 385
rect 40 290 120 300
rect 40 270 50 290
rect 70 280 120 290
rect 70 270 80 280
rect 40 260 80 270
rect 0 220 80 240
rect 60 30 80 220
rect 145 130 165 425
rect 185 185 225 195
rect 185 165 195 185
rect 215 165 225 185
rect 185 155 225 165
rect 145 120 185 130
rect 145 100 155 120
rect 175 100 185 120
rect 145 90 185 100
rect 205 70 225 155
rect 145 50 225 70
rect 145 30 165 50
rect -50 20 -5 30
rect -50 -50 -35 20
rect -15 -50 -5 20
rect -50 -65 -5 -50
rect 60 20 100 30
rect 60 -50 70 20
rect 90 -50 100 20
rect 60 -60 100 -50
rect 125 20 165 30
rect 125 -50 135 20
rect 155 -50 165 20
rect 125 -60 165 -50
rect 190 20 235 30
rect 190 -50 200 20
rect 220 -50 235 20
rect 190 -60 235 -50
rect 20 -110 60 -100
rect 20 -180 30 -110
rect 50 -180 60 -110
rect 20 -190 60 -180
rect 125 -110 165 -100
rect 125 -180 135 -110
rect 155 -180 165 -110
rect 125 -190 165 -180
rect -50 -220 235 -210
rect -50 -230 -15 -220
rect -25 -240 -15 -230
rect 5 -230 90 -220
rect 5 -240 15 -230
rect -25 -245 15 -240
rect 80 -240 90 -230
rect 110 -230 235 -220
rect 110 -240 120 -230
rect 80 -245 120 -240
<< viali >>
rect 30 1285 50 1355
rect 135 1285 155 1355
rect 95 1155 115 1225
rect 95 675 115 745
rect -35 435 -15 505
rect 200 435 220 505
rect -35 -50 -15 20
rect 200 -50 220 20
rect 30 -180 50 -110
rect 135 -180 155 -110
<< metal1 >>
rect -50 1355 235 1370
rect -50 1285 30 1355
rect 50 1285 135 1355
rect 155 1285 235 1355
rect -50 1270 235 1285
rect 85 1225 125 1270
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 745 125 1155
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect -50 20 -5 435
rect -50 -50 -35 20
rect -15 -50 -5 20
rect -50 -95 -5 -50
rect 190 505 235 515
rect 190 435 200 505
rect 220 435 235 505
rect 190 20 235 435
rect 190 -50 200 20
rect 220 -50 235 20
rect 190 -95 235 -50
rect -50 -110 235 -95
rect -50 -180 30 -110
rect 50 -180 135 -110
rect 155 -180 235 -110
rect -50 -195 235 -180
<< labels >>
rlabel locali 235 710 235 710 3 Q
rlabel locali -50 710 -50 710 7 D
rlabel metal1 -50 -150 -50 -150 7 VN
rlabel locali -50 -220 -50 -220 7 CLK
rlabel locali 235 1190 235 1190 3 Qn
rlabel locali -50 1190 -50 1190 7 Dn
rlabel metal1 -50 1325 -50 1325 7 VP
<< end >>
