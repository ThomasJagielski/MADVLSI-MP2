* SPICE3 file created from shift_register_final.ext - technology: sky130A

.subckt inverter A Y VP VN CLK
X0 Y A VP VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=1e+12p ps=6e+06u w=1e+06u l=150000u
X1 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X2 Y A VN VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
.ends

.subckt CSRL_D_FF_width_1 Dn D Qn Q CLK VP VN
X0 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=2e+12p pd=1.2e+07u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X1 Qn Q a_290_2280# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X2 a_30_840# CLK VN VN sky130_fd_pr__nfet_01v8 ad=2.5e+11p pd=2.5e+06u as=0p ps=0u w=1e+06u l=150000u
X3 VP a_30_1320# a_30_2280# VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X4 a_290_1320# CLK VP VP sky130_fd_pr__pfet_01v8 ad=2.5e+11p pd=2.5e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_30_1320# CLK D VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X6 a_30_2280# a_30_1320# a_30_n140# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X7 Qn CLK a_30_2280# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 Q CLK a_30_1320# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X9 a_290_2280# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 Q Qn a_290_1320# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X11 VP a_30_2280# a_30_1320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 a_30_n140# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X13 a_30_2280# CLK Dn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X14 a_30_1320# a_30_2280# a_30_840# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VN Qn Q VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends


* Top level circuit shift_register_final

Xinverter_0 D inverter_0/Y VP VN CLK inverter
XCSRL_D_FF_width_1_0 inverter_0/Y D CSRL_D_FF_width_1_1/Dn CSRL_D_FF_width_1_1/D CLK
+ VP VN CSRL_D_FF_width_1
XCSRL_D_FF_width_1_1 CSRL_D_FF_width_1_1/Dn CSRL_D_FF_width_1_1/D CSRL_D_FF_width_1_2/Dn
+ CSRL_D_FF_width_1_2/D CLK VP VN CSRL_D_FF_width_1
XCSRL_D_FF_width_1_2 CSRL_D_FF_width_1_2/Dn CSRL_D_FF_width_1_2/D CSRL_D_FF_width_1_3/Dn
+ CSRL_D_FF_width_1_3/D CLK VP VN CSRL_D_FF_width_1
XCSRL_D_FF_width_1_3 CSRL_D_FF_width_1_3/Dn CSRL_D_FF_width_1_3/D Qn Q CLK VP VN CSRL_D_FF_width_1
.end

