magic
tech sky130A
timestamp 1614652211
<< nwell >>
rect -70 640 255 1390
<< nmos >>
rect 0 420 15 520
rect 40 420 55 520
rect 105 420 120 520
rect 170 420 185 520
rect 0 -70 15 30
rect 40 -70 55 30
rect 105 -70 120 30
rect 170 -70 185 30
<< pmos >>
rect 0 1140 15 1240
rect 65 1140 80 1240
rect 130 1140 145 1240
rect 170 1140 185 1240
rect 0 660 15 760
rect 65 660 80 760
rect 130 660 145 760
rect 170 660 185 760
<< ndiff >>
rect -50 505 0 520
rect -50 435 -35 505
rect -15 435 0 505
rect -50 420 0 435
rect 15 420 40 520
rect 55 505 105 520
rect 55 435 70 505
rect 90 435 105 505
rect 55 420 105 435
rect 120 505 170 520
rect 120 435 135 505
rect 155 435 170 505
rect 120 420 170 435
rect 185 505 235 520
rect 185 435 200 505
rect 220 435 235 505
rect 185 420 235 435
rect -50 15 0 30
rect -50 -55 -35 15
rect -15 -55 0 15
rect -50 -70 0 -55
rect 15 -70 40 30
rect 55 15 105 30
rect 55 -55 70 15
rect 90 -55 105 15
rect 55 -70 105 -55
rect 120 15 170 30
rect 120 -55 135 15
rect 155 -55 170 15
rect 120 -70 170 -55
rect 185 15 235 30
rect 185 -55 200 15
rect 220 -55 235 15
rect 185 -70 235 -55
<< pdiff >>
rect -50 1225 0 1240
rect -50 1155 -35 1225
rect -15 1155 0 1225
rect -50 1140 0 1155
rect 15 1225 65 1240
rect 15 1155 30 1225
rect 50 1155 65 1225
rect 15 1140 65 1155
rect 80 1225 130 1240
rect 80 1155 95 1225
rect 115 1155 130 1225
rect 80 1140 130 1155
rect 145 1140 170 1240
rect 185 1225 235 1240
rect 185 1155 200 1225
rect 220 1155 235 1225
rect 185 1140 235 1155
rect -50 745 0 760
rect -50 675 -35 745
rect -15 675 0 745
rect -50 660 0 675
rect 15 745 65 760
rect 15 675 30 745
rect 50 675 65 745
rect 15 660 65 675
rect 80 745 130 760
rect 80 675 95 745
rect 115 675 130 745
rect 80 660 130 675
rect 145 660 170 760
rect 185 745 235 760
rect 185 675 200 745
rect 220 675 235 745
rect 185 660 235 675
<< ndiffc >>
rect -35 435 -15 505
rect 70 435 90 505
rect 135 435 155 505
rect 200 435 220 505
rect -35 -55 -15 15
rect 70 -55 90 15
rect 135 -55 155 15
rect 200 -55 220 15
<< pdiffc >>
rect -35 1155 -15 1225
rect 30 1155 50 1225
rect 95 1155 115 1225
rect 200 1155 220 1225
rect -35 675 -15 745
rect 30 675 50 745
rect 95 675 115 745
rect 200 675 220 745
<< psubdiff >>
rect 15 -115 65 -100
rect 15 -185 30 -115
rect 50 -185 65 -115
rect 15 -200 65 -185
rect 120 -115 170 -100
rect 120 -185 135 -115
rect 155 -185 170 -115
rect 120 -200 170 -185
<< nsubdiff >>
rect 15 1355 65 1370
rect 15 1285 30 1355
rect 50 1285 65 1355
rect 15 1270 65 1285
rect 120 1355 170 1370
rect 120 1285 135 1355
rect 155 1285 170 1355
rect 120 1270 170 1285
<< psubdiffcont >>
rect 30 -185 50 -115
rect 135 -185 155 -115
<< nsubdiffcont >>
rect 30 1285 50 1355
rect 135 1285 155 1355
<< poly >>
rect 0 1240 15 1255
rect 65 1240 80 1255
rect 130 1240 145 1255
rect 170 1240 185 1255
rect 0 955 15 1140
rect 65 1085 80 1140
rect 130 1130 145 1140
rect 40 1075 80 1085
rect 40 1055 50 1075
rect 70 1055 80 1075
rect 40 1045 80 1055
rect 105 1115 145 1130
rect 170 1130 185 1140
rect 170 1115 200 1130
rect 40 1010 80 1020
rect 40 990 50 1010
rect 70 990 80 1010
rect 40 980 80 990
rect 0 940 40 955
rect 25 790 40 940
rect 0 775 40 790
rect 0 760 15 775
rect 65 760 80 980
rect 105 785 120 1115
rect 185 915 200 1115
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 105 770 145 785
rect 130 760 145 770
rect 170 760 185 810
rect 0 520 15 660
rect 65 650 80 660
rect 130 650 145 660
rect 40 635 80 650
rect 105 635 145 650
rect 40 520 55 635
rect 105 520 120 635
rect 170 520 185 660
rect 0 235 15 420
rect 40 365 55 420
rect 40 355 80 365
rect 40 335 50 355
rect 70 335 80 355
rect 40 325 80 335
rect 40 290 80 300
rect 40 270 50 290
rect 70 270 80 290
rect 40 260 80 270
rect 0 220 40 235
rect 25 95 40 220
rect 0 80 40 95
rect 0 30 15 80
rect 65 55 80 260
rect 40 40 80 55
rect 40 30 55 40
rect 105 30 120 420
rect 170 190 185 420
rect 170 180 225 190
rect 170 160 195 180
rect 215 160 225 180
rect 170 150 225 160
rect 145 115 185 125
rect 145 95 155 115
rect 175 95 185 115
rect 145 85 185 95
rect 170 30 185 85
rect 0 -215 15 -70
rect 40 -85 55 -70
rect 105 -215 120 -70
rect 170 -85 185 -70
rect -25 -225 15 -215
rect -25 -245 -15 -225
rect 5 -245 15 -225
rect -25 -255 15 -245
rect 80 -225 120 -215
rect 80 -245 90 -225
rect 110 -245 120 -225
rect 80 -255 120 -245
<< polycont >>
rect 50 1055 70 1075
rect 50 990 70 1010
rect 195 885 215 905
rect 155 820 175 840
rect 50 335 70 355
rect 50 270 70 290
rect 195 160 215 180
rect 155 95 175 115
rect -15 -245 5 -225
rect 90 -245 110 -225
<< locali >>
rect 20 1355 60 1365
rect 20 1285 30 1355
rect 50 1285 60 1355
rect 20 1275 60 1285
rect 125 1355 165 1365
rect 125 1285 135 1355
rect 155 1285 165 1355
rect 125 1275 165 1285
rect -50 1225 -5 1235
rect -50 1155 -35 1225
rect -15 1155 -5 1225
rect -50 1145 -5 1155
rect 20 1225 60 1235
rect 20 1155 30 1225
rect 50 1155 60 1225
rect 20 1145 60 1155
rect 85 1225 125 1235
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 1145 125 1155
rect 190 1225 235 1235
rect 190 1155 200 1225
rect 220 1155 235 1225
rect 190 1145 235 1155
rect 40 1125 60 1145
rect 190 1125 210 1145
rect 40 1105 120 1125
rect 40 1075 80 1085
rect 40 1065 50 1075
rect 0 1055 50 1065
rect 70 1055 80 1075
rect 0 1045 80 1055
rect 0 960 20 1045
rect 100 1020 120 1105
rect 40 1010 120 1020
rect 40 990 50 1010
rect 70 1000 120 1010
rect 145 1105 210 1125
rect 70 990 80 1000
rect 40 980 80 990
rect 0 940 40 960
rect 20 755 40 940
rect 145 850 165 1105
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 205 755 225 875
rect -50 745 -5 755
rect -50 675 -35 745
rect -15 675 -5 745
rect -50 665 -5 675
rect 20 745 60 755
rect 20 675 30 745
rect 50 675 60 745
rect 20 665 60 675
rect 85 745 125 755
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect 190 745 235 755
rect 190 675 200 745
rect 220 675 235 745
rect 190 665 235 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect 40 515 60 665
rect 190 640 210 665
rect 145 620 210 640
rect 145 515 165 620
rect 40 505 100 515
rect 40 495 70 505
rect -50 425 -5 435
rect 60 435 70 495
rect 90 435 100 505
rect 60 425 100 435
rect 125 505 165 515
rect 125 435 135 505
rect 155 435 165 505
rect 125 425 165 435
rect 190 505 235 515
rect 190 435 200 505
rect 220 435 235 505
rect 190 425 235 435
rect 80 405 100 425
rect 80 385 120 405
rect 40 355 80 365
rect 40 345 50 355
rect 0 335 50 345
rect 70 335 80 355
rect 0 325 80 335
rect 0 240 20 325
rect 100 300 120 385
rect 40 290 120 300
rect 40 270 50 290
rect 70 280 120 290
rect 70 270 80 280
rect 40 260 80 270
rect 0 220 80 240
rect 60 25 80 220
rect 145 125 165 425
rect 185 180 225 190
rect 185 160 195 180
rect 215 160 225 180
rect 185 150 225 160
rect 145 115 185 125
rect 145 95 155 115
rect 175 95 185 115
rect 145 85 185 95
rect 205 65 225 150
rect 145 45 225 65
rect 145 25 165 45
rect -50 15 -5 25
rect -50 -55 -35 15
rect -15 -55 -5 15
rect -50 -70 -5 -55
rect 60 15 100 25
rect 60 -55 70 15
rect 90 -55 100 15
rect 60 -65 100 -55
rect 125 15 165 25
rect 125 -55 135 15
rect 155 -55 165 15
rect 125 -65 165 -55
rect 190 15 235 25
rect 190 -55 200 15
rect 220 -55 235 15
rect 190 -65 235 -55
rect 20 -115 60 -105
rect 20 -185 30 -115
rect 50 -185 60 -115
rect 20 -195 60 -185
rect 125 -115 165 -105
rect 125 -185 135 -115
rect 155 -185 165 -115
rect 125 -195 165 -185
rect -50 -225 235 -215
rect -50 -235 -15 -225
rect -25 -245 -15 -235
rect 5 -235 90 -225
rect 5 -245 15 -235
rect -25 -255 15 -245
rect 80 -245 90 -235
rect 110 -235 235 -225
rect 110 -245 120 -235
rect 80 -255 120 -245
<< viali >>
rect 30 1285 50 1355
rect 135 1285 155 1355
rect 95 1155 115 1225
rect 95 675 115 745
rect -35 435 -15 505
rect 200 435 220 505
rect -35 -55 -15 15
rect 200 -55 220 15
rect 30 -185 50 -115
rect 135 -185 155 -115
<< metal1 >>
rect -50 1355 235 1370
rect -50 1285 30 1355
rect 50 1285 135 1355
rect 155 1285 235 1355
rect -50 1270 235 1285
rect 85 1225 125 1270
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 745 125 1155
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect -50 15 -5 435
rect -50 -55 -35 15
rect -15 -55 -5 15
rect -50 -100 -5 -55
rect 190 505 235 515
rect 190 435 200 505
rect 220 435 235 505
rect 190 15 235 435
rect 190 -55 200 15
rect 220 -55 235 15
rect 190 -100 235 -55
rect -50 -115 235 -100
rect -50 -185 30 -115
rect 50 -185 135 -115
rect 155 -185 235 -115
rect -50 -200 235 -185
<< labels >>
rlabel locali 235 710 235 710 3 Q
rlabel locali -50 710 -50 710 7 D
rlabel locali 235 1190 235 1190 3 Qn
rlabel locali -50 1190 -50 1190 7 Dn
rlabel metal1 -50 1325 -50 1325 7 VP
rlabel metal1 -50 -155 -50 -155 7 VN
rlabel locali -50 -225 -50 -225 7 CLK
<< end >>
