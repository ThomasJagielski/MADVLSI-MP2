magic
tech sky130A
timestamp 1614621003
<< nwell >>
rect -70 655 85 1240
<< nmos >>
rect 0 230 15 330
<< pmos >>
rect 0 890 15 1090
<< ndiff >>
rect -50 315 0 330
rect -50 245 -35 315
rect -15 245 0 315
rect -50 230 0 245
rect 15 315 65 330
rect 15 245 30 315
rect 50 245 65 315
rect 15 230 65 245
<< pdiff >>
rect -50 1075 0 1090
rect -50 1005 -35 1075
rect -15 1005 0 1075
rect -50 975 0 1005
rect -50 905 -35 975
rect -15 905 0 975
rect -50 890 0 905
rect 15 1075 65 1090
rect 15 1005 30 1075
rect 50 1005 65 1075
rect 15 975 65 1005
rect 15 905 30 975
rect 50 905 65 975
rect 15 890 65 905
<< ndiffc >>
rect -35 245 -15 315
rect 30 245 50 315
<< pdiffc >>
rect -35 1005 -15 1075
rect -35 905 -15 975
rect 30 1005 50 1075
rect 30 905 50 975
<< psubdiff >>
rect -50 -45 0 -30
rect -50 -115 -35 -45
rect -15 -115 0 -45
rect -50 -130 0 -115
<< nsubdiff >>
rect -50 1205 0 1220
rect -50 1135 -35 1205
rect -15 1135 0 1205
rect -50 1120 0 1135
<< psubdiffcont >>
rect -35 -115 -15 -45
<< nsubdiffcont >>
rect -35 1135 -15 1205
<< poly >>
rect 0 1090 15 1105
rect 0 875 15 890
rect -45 865 15 875
rect -45 845 -35 865
rect -15 860 15 865
rect -15 845 -5 860
rect -45 835 -5 845
rect -45 620 -30 835
rect -45 610 35 620
rect -45 605 5 610
rect -45 355 -30 605
rect -5 590 5 605
rect 25 590 35 610
rect -5 580 35 590
rect -45 340 15 355
rect 0 330 15 340
rect 0 215 15 230
<< polycont >>
rect -35 845 -15 865
rect 5 590 25 610
<< locali >>
rect -45 1205 -5 1215
rect -45 1135 -35 1205
rect -15 1135 -5 1205
rect -45 1125 -5 1135
rect -45 1075 -5 1085
rect -45 1005 -35 1075
rect -15 1005 -5 1075
rect -45 975 -5 1005
rect -45 905 -35 975
rect -15 905 -5 975
rect -45 895 -5 905
rect 20 1075 65 1085
rect 20 1005 30 1075
rect 50 1005 65 1075
rect 20 995 65 1005
rect 20 975 60 995
rect 20 905 30 975
rect 50 905 60 975
rect 20 900 60 905
rect -45 865 -5 875
rect -45 845 -35 865
rect -15 845 -5 865
rect -45 835 -5 845
rect -45 770 -25 835
rect 20 815 40 900
rect -50 680 -25 770
rect -5 795 40 815
rect -5 660 15 795
rect -45 640 15 660
rect 35 680 65 770
rect -45 560 -25 640
rect 35 620 55 680
rect -5 610 55 620
rect -5 590 5 610
rect 25 600 55 610
rect 25 590 35 600
rect -5 580 35 590
rect -45 540 40 560
rect 20 325 40 540
rect -45 315 -5 325
rect -45 245 -35 315
rect -15 245 -5 315
rect -45 235 -5 245
rect 20 315 60 325
rect 20 245 30 315
rect 50 245 60 315
rect 20 235 60 245
rect -45 -45 -5 -35
rect -45 -115 -35 -45
rect -15 -115 -5 -45
rect -45 -125 -5 -115
rect -50 -165 65 -145
<< viali >>
rect -35 1135 -15 1205
rect -35 1005 -15 1075
rect -35 905 -15 975
rect -35 245 -15 315
rect -35 -115 -15 -45
<< metal1 >>
rect -50 1205 65 1220
rect -50 1135 -35 1205
rect -15 1135 65 1205
rect -50 1120 65 1135
rect -45 1075 -5 1120
rect -45 1005 -35 1075
rect -15 1005 -5 1075
rect -45 975 -5 1005
rect -45 905 -35 975
rect -15 905 -5 975
rect -45 895 -5 905
rect -45 315 -5 325
rect -45 245 -35 315
rect -15 245 -5 315
rect -45 -30 -5 245
rect -50 -45 65 -30
rect -50 -115 -35 -45
rect -15 -115 65 -45
rect -50 -130 65 -115
<< labels >>
rlabel metal1 -50 1170 -50 1170 7 VP
port 3 w
rlabel locali -50 725 -50 725 7 A
port 1 w
rlabel locali 65 1040 65 1040 3 Y
port 2 e
rlabel metal1 -50 -80 -50 -80 7 VN
port 4 w
rlabel locali -50 -155 -50 -155 7 CLK
port 5 w
rlabel locali 65 725 65 725 3 Ao
port 6 e
<< end >>
