magic
tech sky130A
timestamp 1614625195
<< nwell >>
rect -70 705 85 1455
<< nmos >>
rect 0 230 15 330
<< pmos >>
rect 0 1105 15 1305
<< ndiff >>
rect -50 315 0 330
rect -50 245 -35 315
rect -15 245 0 315
rect -50 230 0 245
rect 15 315 65 330
rect 15 245 30 315
rect 50 245 65 315
rect 15 230 65 245
<< pdiff >>
rect -50 1290 0 1305
rect -50 1220 -35 1290
rect -15 1220 0 1290
rect -50 1190 0 1220
rect -50 1120 -35 1190
rect -15 1120 0 1190
rect -50 1105 0 1120
rect 15 1290 65 1305
rect 15 1220 30 1290
rect 50 1220 65 1290
rect 15 1190 65 1220
rect 15 1120 30 1190
rect 50 1120 65 1190
rect 15 1105 65 1120
<< ndiffc >>
rect -35 245 -15 315
rect 30 245 50 315
<< pdiffc >>
rect -35 1220 -15 1290
rect -35 1120 -15 1190
rect 30 1220 50 1290
rect 30 1120 50 1190
<< psubdiff >>
rect -50 -45 0 -30
rect -50 -115 -35 -45
rect -15 -115 0 -45
rect -50 -130 0 -115
<< nsubdiff >>
rect -50 1420 0 1435
rect -50 1350 -35 1420
rect -15 1350 0 1420
rect -50 1335 0 1350
<< psubdiffcont >>
rect -35 -115 -15 -45
<< nsubdiffcont >>
rect -35 1350 -15 1420
<< poly >>
rect 0 1305 15 1320
rect 0 1090 15 1105
rect -45 1080 15 1090
rect -45 1060 -35 1080
rect -15 1075 15 1080
rect -15 1060 -5 1075
rect -45 1050 -5 1060
rect -45 670 -30 1050
rect -45 660 35 670
rect -45 655 5 660
rect -45 355 -30 655
rect -5 640 5 655
rect 25 640 35 660
rect -5 630 35 640
rect -45 340 15 355
rect 0 330 15 340
rect 0 215 15 230
<< polycont >>
rect -35 1060 -15 1080
rect 5 640 25 660
<< locali >>
rect -45 1420 -5 1430
rect -45 1350 -35 1420
rect -15 1350 -5 1420
rect -45 1340 -5 1350
rect -45 1290 -5 1300
rect -45 1220 -35 1290
rect -15 1220 -5 1290
rect -45 1190 -5 1220
rect -45 1120 -35 1190
rect -15 1120 -5 1190
rect -45 1110 -5 1120
rect 20 1290 65 1300
rect 20 1220 30 1290
rect 50 1220 65 1290
rect 20 1210 65 1220
rect 20 1190 60 1210
rect 20 1120 30 1190
rect 50 1120 60 1190
rect 20 1115 60 1120
rect -45 1080 -5 1090
rect -45 1060 -35 1080
rect -15 1060 -5 1080
rect -45 1050 -5 1060
rect -45 820 -25 1050
rect 20 1030 40 1115
rect -50 730 -25 820
rect -5 1010 40 1030
rect -5 710 15 1010
rect -45 690 15 710
rect 35 730 65 820
rect -45 365 -25 690
rect 35 670 55 730
rect -5 660 55 670
rect -5 640 5 660
rect 25 650 55 660
rect 25 640 35 650
rect -5 630 35 640
rect -45 345 40 365
rect 20 325 40 345
rect -45 315 -5 325
rect -45 245 -35 315
rect -15 245 -5 315
rect -45 235 -5 245
rect 20 315 60 325
rect 20 245 30 315
rect 50 245 60 315
rect 20 235 60 245
rect -45 -45 -5 -35
rect -45 -115 -35 -45
rect -15 -115 -5 -45
rect -45 -125 -5 -115
rect -50 -165 65 -145
<< viali >>
rect -35 1350 -15 1420
rect -35 1220 -15 1290
rect -35 1120 -15 1190
rect -35 245 -15 315
rect -35 -115 -15 -45
<< metal1 >>
rect -50 1420 65 1435
rect -50 1350 -35 1420
rect -15 1350 65 1420
rect -50 1335 65 1350
rect -45 1290 -5 1335
rect -45 1220 -35 1290
rect -15 1220 -5 1290
rect -45 1190 -5 1220
rect -45 1120 -35 1190
rect -15 1120 -5 1190
rect -45 1110 -5 1120
rect -45 315 -5 325
rect -45 245 -35 315
rect -15 245 -5 315
rect -45 -30 -5 245
rect -50 -45 65 -30
rect -50 -115 -35 -45
rect -15 -115 65 -45
rect -50 -130 65 -115
<< labels >>
rlabel metal1 -50 -80 -50 -80 7 VN
port 4 w
rlabel locali -50 -155 -50 -155 7 CLK
port 5 w
rlabel metal1 -50 1385 -50 1385 7 VP
port 3 w
rlabel locali 65 1255 65 1255 3 Y
port 2 e
rlabel locali -50 775 -50 775 7 A
port 1 w
rlabel locali 65 775 65 775 3 Ao
port 6 e
<< end >>
