magic
tech sky130A
timestamp 1614619059
<< nwell >>
rect -70 640 255 1225
<< nmos >>
rect 0 355 15 555
rect 40 355 55 555
rect 105 455 120 555
rect 170 455 185 555
rect 0 -15 15 185
rect 40 -15 55 185
rect 105 -15 120 85
rect 170 -15 185 85
<< pmos >>
rect 0 975 15 1075
rect 65 975 80 1075
rect 130 975 145 1075
rect 170 975 185 1075
rect 0 660 15 760
rect 65 660 80 760
rect 130 660 145 760
rect 170 660 185 760
<< ndiff >>
rect -50 540 0 555
rect -50 470 -35 540
rect -15 470 0 540
rect -50 440 0 470
rect -50 370 -35 440
rect -15 370 0 440
rect -50 355 0 370
rect 15 355 40 555
rect 55 540 105 555
rect 55 470 70 540
rect 90 470 105 540
rect 55 455 105 470
rect 120 540 170 555
rect 120 470 135 540
rect 155 470 170 540
rect 120 455 170 470
rect 185 540 235 555
rect 185 470 200 540
rect 220 470 235 540
rect 185 455 235 470
rect 55 355 80 455
rect -50 170 0 185
rect -50 100 -35 170
rect -15 100 0 170
rect -50 70 0 100
rect -50 0 -35 70
rect -15 0 0 70
rect -50 -15 0 0
rect 15 -15 40 185
rect 55 85 80 185
rect 55 70 105 85
rect 55 0 70 70
rect 90 0 105 70
rect 55 -15 105 0
rect 120 70 170 85
rect 120 0 135 70
rect 155 0 170 70
rect 120 -15 170 0
rect 185 70 235 85
rect 185 0 200 70
rect 220 0 235 70
rect 185 -15 235 0
<< pdiff >>
rect -50 1060 0 1075
rect -50 990 -35 1060
rect -15 990 0 1060
rect -50 975 0 990
rect 15 1060 65 1075
rect 15 990 30 1060
rect 50 990 65 1060
rect 15 975 65 990
rect 80 1060 130 1075
rect 80 990 95 1060
rect 115 990 130 1060
rect 80 975 130 990
rect 145 975 170 1075
rect 185 1060 235 1075
rect 185 990 200 1060
rect 220 990 235 1060
rect 185 975 235 990
rect -50 745 0 760
rect -50 675 -35 745
rect -15 675 0 745
rect -50 660 0 675
rect 15 745 65 760
rect 15 675 30 745
rect 50 675 65 745
rect 15 660 65 675
rect 80 745 130 760
rect 80 675 95 745
rect 115 675 130 745
rect 80 660 130 675
rect 145 660 170 760
rect 185 745 235 760
rect 185 675 200 745
rect 220 675 235 745
rect 185 660 235 675
<< ndiffc >>
rect -35 470 -15 540
rect -35 370 -15 440
rect 70 470 90 540
rect 135 470 155 540
rect 200 470 220 540
rect -35 100 -15 170
rect -35 0 -15 70
rect 70 0 90 70
rect 135 0 155 70
rect 200 0 220 70
<< pdiffc >>
rect -35 990 -15 1060
rect 30 990 50 1060
rect 95 990 115 1060
rect 200 990 220 1060
rect -35 675 -15 745
rect 30 675 50 745
rect 95 675 115 745
rect 200 675 220 745
<< psubdiff >>
rect 15 -60 65 -45
rect 15 -130 30 -60
rect 50 -130 65 -60
rect 15 -145 65 -130
rect 120 -60 170 -45
rect 120 -130 135 -60
rect 155 -130 170 -60
rect 120 -145 170 -130
<< nsubdiff >>
rect 15 1190 65 1205
rect 15 1120 30 1190
rect 50 1120 65 1190
rect 15 1105 65 1120
rect 120 1190 170 1205
rect 120 1120 135 1190
rect 155 1120 170 1190
rect 120 1105 170 1120
<< psubdiffcont >>
rect 30 -130 50 -60
rect 135 -130 155 -60
<< nsubdiffcont >>
rect 30 1120 50 1190
rect 135 1120 155 1190
<< poly >>
rect 0 1075 15 1090
rect 65 1075 80 1090
rect 130 1075 145 1090
rect 170 1075 185 1090
rect 0 760 15 975
rect 65 920 80 975
rect 130 965 145 975
rect 40 910 80 920
rect 40 890 50 910
rect 70 890 80 910
rect 40 880 80 890
rect 105 950 145 965
rect 40 845 80 855
rect 40 825 50 845
rect 70 825 80 845
rect 40 815 80 825
rect 65 760 80 815
rect 105 785 120 950
rect 170 920 185 975
rect 145 910 185 920
rect 145 890 155 910
rect 175 890 185 910
rect 145 880 185 890
rect 170 845 225 855
rect 170 825 195 845
rect 215 825 225 845
rect 170 815 225 825
rect 105 770 145 785
rect 130 760 145 770
rect 170 760 185 815
rect 0 555 15 660
rect 65 650 80 660
rect 130 650 145 660
rect 40 635 80 650
rect 105 635 145 650
rect 40 555 55 635
rect 105 555 120 635
rect 170 555 185 660
rect 0 185 15 355
rect 40 345 55 355
rect 40 335 80 345
rect 40 315 50 335
rect 70 315 80 335
rect 40 305 80 315
rect 40 270 80 280
rect 40 250 50 270
rect 70 250 80 270
rect 40 240 80 250
rect 40 185 55 240
rect 105 85 120 455
rect 170 430 185 455
rect 145 415 185 430
rect 145 185 160 415
rect 185 240 225 250
rect 185 220 195 240
rect 215 220 225 240
rect 185 210 225 220
rect 145 175 185 185
rect 145 155 155 175
rect 175 155 185 175
rect 145 145 185 155
rect 210 120 225 210
rect 170 105 225 120
rect 170 85 185 105
rect 0 -160 15 -15
rect 40 -30 55 -15
rect 105 -160 120 -15
rect 170 -30 185 -15
rect -25 -170 15 -160
rect -25 -190 -15 -170
rect 5 -190 15 -170
rect -25 -200 15 -190
rect 80 -170 120 -160
rect 80 -190 90 -170
rect 110 -190 120 -170
rect 80 -200 120 -190
<< polycont >>
rect 50 890 70 910
rect 50 825 70 845
rect 155 890 175 910
rect 195 825 215 845
rect 50 315 70 335
rect 50 250 70 270
rect 195 220 215 240
rect 155 155 175 175
rect -15 -190 5 -170
rect 90 -190 110 -170
<< locali >>
rect 20 1190 60 1200
rect 20 1120 30 1190
rect 50 1120 60 1190
rect 20 1110 60 1120
rect 125 1190 165 1200
rect 125 1120 135 1190
rect 155 1120 165 1190
rect 125 1110 165 1120
rect -50 1060 -5 1070
rect -50 990 -35 1060
rect -15 990 -5 1060
rect -50 980 -5 990
rect 20 1060 60 1070
rect 20 990 30 1060
rect 50 990 60 1060
rect 20 980 60 990
rect 85 1060 125 1070
rect 85 990 95 1060
rect 115 990 125 1060
rect 85 980 125 990
rect 190 1060 235 1070
rect 190 990 200 1060
rect 220 990 235 1060
rect 190 980 235 990
rect 40 960 60 980
rect 40 940 120 960
rect 40 910 80 920
rect 40 900 50 910
rect 0 890 50 900
rect 70 890 80 910
rect 0 880 80 890
rect 0 795 20 880
rect 100 855 120 940
rect 40 845 120 855
rect 40 825 50 845
rect 70 835 120 845
rect 145 910 185 920
rect 145 890 155 910
rect 175 890 185 910
rect 145 880 185 890
rect 70 825 80 835
rect 40 815 80 825
rect 0 775 40 795
rect 20 755 40 775
rect 145 755 165 880
rect 205 855 225 980
rect 185 845 225 855
rect 185 825 195 845
rect 215 825 225 845
rect 185 815 225 825
rect -50 745 -5 755
rect -50 675 -35 745
rect -15 675 -5 745
rect -50 665 -5 675
rect 20 745 60 755
rect 20 675 30 745
rect 50 675 60 745
rect 20 665 60 675
rect 85 745 125 755
rect 85 675 95 745
rect 115 675 125 745
rect 145 745 235 755
rect 145 735 200 745
rect 85 665 125 675
rect 190 675 200 735
rect 220 675 235 745
rect 190 665 235 675
rect 40 550 60 665
rect 190 640 210 665
rect 145 620 210 640
rect 145 550 165 620
rect -50 540 -5 550
rect -50 470 -35 540
rect -15 470 -5 540
rect 40 540 100 550
rect 40 530 70 540
rect -50 440 -5 470
rect 60 470 70 530
rect 90 470 100 540
rect 60 460 100 470
rect 125 540 165 550
rect 125 470 135 540
rect 155 470 165 540
rect 125 460 165 470
rect 190 540 235 550
rect 190 470 200 540
rect 220 470 235 540
rect 190 460 235 470
rect -50 370 -35 440
rect -15 370 -5 440
rect -50 360 -5 370
rect 80 385 100 460
rect 80 365 120 385
rect 40 335 80 345
rect 40 325 50 335
rect 0 315 50 325
rect 70 315 80 335
rect 0 305 80 315
rect 0 220 20 305
rect 100 280 120 365
rect 40 270 120 280
rect 40 250 50 270
rect 70 260 120 270
rect 70 250 80 260
rect 40 240 80 250
rect 140 250 160 460
rect 140 240 225 250
rect 140 230 195 240
rect 185 220 195 230
rect 215 220 225 240
rect 0 200 35 220
rect 185 210 225 220
rect -50 170 -5 180
rect -50 100 -35 170
rect -15 100 -5 170
rect -50 70 -5 100
rect -50 0 -35 70
rect -15 0 -5 70
rect 15 80 35 200
rect 145 175 185 185
rect 145 155 155 175
rect 175 155 185 175
rect 145 145 185 155
rect 145 80 165 145
rect 15 70 100 80
rect 15 60 70 70
rect -50 -10 -5 0
rect 60 0 70 60
rect 90 0 100 70
rect 60 -10 100 0
rect 125 70 165 80
rect 125 0 135 70
rect 155 0 165 70
rect 125 -10 165 0
rect 190 70 235 80
rect 190 0 200 70
rect 220 0 235 70
rect 190 -10 235 0
rect 20 -60 60 -50
rect 20 -130 30 -60
rect 50 -130 60 -60
rect 20 -140 60 -130
rect 125 -60 165 -50
rect 125 -130 135 -60
rect 155 -130 165 -60
rect 125 -140 165 -130
rect -50 -170 235 -160
rect -50 -180 -15 -170
rect -25 -190 -15 -180
rect 5 -180 90 -170
rect 5 -190 15 -180
rect -25 -200 15 -190
rect 80 -190 90 -180
rect 110 -180 235 -170
rect 110 -190 120 -180
rect 80 -200 120 -190
<< viali >>
rect 30 1120 50 1190
rect 135 1120 155 1190
rect 95 990 115 1060
rect 95 675 115 745
rect -35 470 -15 540
rect 200 470 220 540
rect -35 370 -15 440
rect -35 100 -15 170
rect -35 0 -15 70
rect 200 0 220 70
rect 30 -130 50 -60
rect 135 -130 155 -60
<< metal1 >>
rect -50 1190 235 1205
rect -50 1120 30 1190
rect 50 1120 135 1190
rect 155 1120 235 1190
rect -50 1105 235 1120
rect 85 1060 125 1105
rect 85 990 95 1060
rect 115 990 125 1060
rect 85 745 125 990
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect -50 540 -5 550
rect -50 470 -35 540
rect -15 470 -5 540
rect -50 440 -5 470
rect -50 370 -35 440
rect -15 370 -5 440
rect -50 170 -5 370
rect -50 100 -35 170
rect -15 100 -5 170
rect -50 70 -5 100
rect -50 0 -35 70
rect -15 0 -5 70
rect -50 -45 -5 0
rect 190 540 235 550
rect 190 470 200 540
rect 220 470 235 540
rect 190 70 235 470
rect 190 0 200 70
rect 220 0 235 70
rect 190 -45 235 0
rect -50 -60 235 -45
rect -50 -130 30 -60
rect 50 -130 135 -60
rect 155 -130 235 -60
rect -50 -145 235 -130
<< labels >>
rlabel locali 235 1025 235 1025 3 Qn
rlabel locali 235 710 235 710 3 Q
rlabel locali -50 710 -50 710 7 D
rlabel locali -50 1025 -50 1025 7 Dn
rlabel metal1 -50 1160 -50 1160 7 VP
rlabel locali -50 -170 -50 -170 7 CLK
rlabel metal1 -50 -100 -50 -100 7 VN
<< end >>
