magic
tech sky130A
timestamp 1614628828
<< locali >>
rect 1135 1385 1150 1475
rect 55 905 80 995
rect 1135 905 1150 995
rect 55 10 70 30
<< metal1 >>
rect 55 1510 70 1610
rect 55 45 70 145
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_3
timestamp 1614455318
transform 1 0 915 0 1 240
box -70 -245 255 1395
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_2
timestamp 1614455318
transform 1 0 680 0 1 240
box -70 -245 255 1395
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_1
timestamp 1614455318
transform 1 0 445 0 1 240
box -70 -245 255 1395
use inverter  inverter_0
timestamp 1614625195
transform 1 0 105 0 1 175
box -70 -165 85 1455
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_0
timestamp 1614455318
transform 1 0 210 0 1 240
box -70 -245 255 1395
<< labels >>
rlabel locali 55 950 55 950 7 D
rlabel metal1 55 1560 55 1560 7 VP
rlabel metal1 55 95 55 95 7 VN
rlabel locali 55 20 55 20 7 CLK
rlabel locali 1150 950 1150 950 3 Q
rlabel locali 1150 1430 1150 1430 3 Qn
<< end >>
