magic
tech sky130A
timestamp 1614455710
<< locali >>
rect 20 1390 35 1480
rect 995 1390 1010 1480
rect 20 910 35 1000
rect 995 910 1010 1000
rect 20 15 35 35
<< metal1 >>
rect 20 1515 50 1615
rect 20 50 50 150
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_3 ~/Documents/MADVLSI-MP2/layout/width_1_transistors
timestamp 1614455318
transform 1 0 775 0 1 245
box -70 -245 255 1395
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_2
timestamp 1614455318
transform 1 0 540 0 1 245
box -70 -245 255 1395
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_1
timestamp 1614455318
transform 1 0 305 0 1 245
box -70 -245 255 1395
use CSRL_D_FF_width_1  CSRL_D_FF_width_1_0
timestamp 1614455318
transform 1 0 70 0 1 245
box -70 -245 255 1395
<< labels >>
rlabel metal1 20 1565 20 1565 7 VP
rlabel locali 20 1435 20 1435 7 Dn
rlabel locali 20 955 20 955 7 D
rlabel metal1 20 100 20 100 7 VN
rlabel locali 20 25 20 25 7 CLK
rlabel locali 1010 955 1010 955 3 Q
rlabel locali 1010 1435 1010 1435 3 Qn
<< end >>
