magic
tech sky130A
timestamp 1614281118
<< nwell >>
rect -70 640 255 1380
<< nmos >>
rect 0 320 15 520
rect 40 320 55 520
rect 105 320 120 420
rect 170 320 185 420
rect 0 -115 15 85
rect 40 -115 55 85
rect 105 -15 120 85
rect 170 -15 185 85
<< pmos >>
rect 0 1125 15 1225
rect 65 1125 80 1225
rect 130 1125 145 1225
rect 170 1125 185 1225
rect 0 660 15 760
rect 65 660 80 760
rect 130 660 145 760
rect 170 660 185 760
<< ndiff >>
rect -50 505 0 520
rect -50 435 -35 505
rect -15 435 0 505
rect -50 405 0 435
rect -50 335 -35 405
rect -15 335 0 405
rect -50 320 0 335
rect 15 320 40 520
rect 55 420 80 520
rect 55 405 105 420
rect 55 335 70 405
rect 90 335 105 405
rect 55 320 105 335
rect 120 405 170 420
rect 120 335 135 405
rect 155 335 170 405
rect 120 320 170 335
rect 185 405 235 420
rect 185 335 200 405
rect 220 335 235 405
rect 185 320 235 335
rect -50 70 0 85
rect -50 0 -35 70
rect -15 0 0 70
rect -50 -30 0 0
rect -50 -100 -35 -30
rect -15 -100 0 -30
rect -50 -115 0 -100
rect 15 -115 40 85
rect 55 70 105 85
rect 55 0 70 70
rect 90 0 105 70
rect 55 -15 105 0
rect 120 70 170 85
rect 120 0 135 70
rect 155 0 170 70
rect 120 -15 170 0
rect 185 70 235 85
rect 185 0 200 70
rect 220 0 235 70
rect 185 -15 235 0
rect 55 -115 80 -15
<< pdiff >>
rect -50 1210 0 1225
rect -50 1140 -35 1210
rect -15 1140 0 1210
rect -50 1125 0 1140
rect 15 1210 65 1225
rect 15 1140 30 1210
rect 50 1140 65 1210
rect 15 1125 65 1140
rect 80 1210 130 1225
rect 80 1140 95 1210
rect 115 1140 130 1210
rect 80 1125 130 1140
rect 145 1125 170 1225
rect 185 1210 235 1225
rect 185 1140 200 1210
rect 220 1140 235 1210
rect 185 1125 235 1140
rect -50 745 0 760
rect -50 675 -35 745
rect -15 675 0 745
rect -50 660 0 675
rect 15 745 65 760
rect 15 675 30 745
rect 50 675 65 745
rect 15 660 65 675
rect 80 745 130 760
rect 80 675 95 745
rect 115 675 130 745
rect 80 660 130 675
rect 145 660 170 760
rect 185 745 235 760
rect 185 675 200 745
rect 220 675 235 745
rect 185 660 235 675
<< ndiffc >>
rect -35 435 -15 505
rect -35 335 -15 405
rect 70 335 90 405
rect 135 335 155 405
rect 200 335 220 405
rect -35 0 -15 70
rect -35 -100 -15 -30
rect 70 0 90 70
rect 135 0 155 70
rect 200 0 220 70
<< pdiffc >>
rect -35 1140 -15 1210
rect 30 1140 50 1210
rect 95 1140 115 1210
rect 200 1140 220 1210
rect -35 675 -15 745
rect 30 675 50 745
rect 95 675 115 745
rect 200 675 220 745
<< psubdiff >>
rect 15 -160 65 -145
rect 15 -230 30 -160
rect 50 -230 65 -160
rect 15 -245 65 -230
rect 120 -160 170 -145
rect 120 -230 135 -160
rect 155 -230 170 -160
rect 120 -245 170 -230
<< nsubdiff >>
rect 15 1340 65 1355
rect 15 1270 30 1340
rect 50 1270 65 1340
rect 15 1255 65 1270
rect 120 1340 170 1355
rect 120 1270 135 1340
rect 155 1270 170 1340
rect 120 1255 170 1270
<< psubdiffcont >>
rect 30 -230 50 -160
rect 135 -230 155 -160
<< nsubdiffcont >>
rect 30 1270 50 1340
rect 135 1270 155 1340
<< poly >>
rect 0 1225 15 1240
rect 65 1225 80 1240
rect 130 1225 145 1240
rect 170 1225 185 1240
rect 0 760 15 1125
rect 65 1070 80 1125
rect 130 1115 145 1125
rect 40 1060 80 1070
rect 40 1040 50 1060
rect 70 1040 80 1060
rect 40 1030 80 1040
rect 105 1100 145 1115
rect 170 1115 185 1125
rect 170 1100 200 1115
rect 40 995 80 1005
rect 40 975 50 995
rect 70 975 80 995
rect 40 965 80 975
rect 65 760 80 965
rect 105 785 120 1100
rect 185 915 200 1100
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 105 770 145 785
rect 130 760 145 770
rect 170 760 185 810
rect 0 520 15 660
rect 65 650 80 660
rect 130 650 145 660
rect 40 635 80 650
rect 105 635 145 650
rect 40 520 55 635
rect 105 420 120 635
rect 170 420 185 660
rect 0 85 15 320
rect 40 250 55 320
rect 40 240 80 250
rect 40 220 50 240
rect 70 220 80 240
rect 40 210 80 220
rect 40 175 80 185
rect 40 155 50 175
rect 70 155 80 175
rect 40 145 80 155
rect 40 85 55 145
rect 105 85 120 320
rect 170 295 185 320
rect 145 280 185 295
rect 145 185 160 280
rect 185 245 225 255
rect 185 225 195 245
rect 215 225 225 245
rect 185 215 225 225
rect 145 175 185 185
rect 145 155 155 175
rect 175 155 185 175
rect 145 145 185 155
rect 210 120 225 215
rect 170 105 225 120
rect 170 85 185 105
rect 0 -260 15 -115
rect 40 -130 55 -115
rect 105 -260 120 -15
rect 170 -30 185 -15
rect -25 -270 15 -260
rect -25 -290 -15 -270
rect 5 -290 15 -270
rect -25 -295 15 -290
rect 80 -270 120 -260
rect 80 -290 90 -270
rect 110 -290 120 -270
rect 80 -295 120 -290
<< polycont >>
rect 50 1040 70 1060
rect 50 975 70 995
rect 195 885 215 905
rect 155 820 175 840
rect 50 220 70 240
rect 50 155 70 175
rect 195 225 215 245
rect 155 155 175 175
rect -15 -290 5 -270
rect 90 -290 110 -270
<< locali >>
rect 20 1340 60 1350
rect 20 1270 30 1340
rect 50 1270 60 1340
rect 20 1260 60 1270
rect 125 1340 165 1350
rect 125 1270 135 1340
rect 155 1270 165 1340
rect 125 1260 165 1270
rect -50 1210 -5 1220
rect -50 1140 -35 1210
rect -15 1140 -5 1210
rect -50 1130 -5 1140
rect 20 1210 60 1220
rect 20 1140 30 1210
rect 50 1140 60 1210
rect 20 1130 60 1140
rect 85 1210 125 1220
rect 85 1140 95 1210
rect 115 1140 125 1210
rect 85 1130 125 1140
rect 190 1210 235 1220
rect 190 1140 200 1210
rect 220 1140 235 1210
rect 190 1130 235 1140
rect 40 1110 60 1130
rect 190 1110 210 1130
rect 40 1090 120 1110
rect 40 1060 80 1070
rect 40 1050 50 1060
rect 0 1040 50 1050
rect 70 1040 80 1060
rect 0 1030 80 1040
rect 0 945 20 1030
rect 100 1005 120 1090
rect 40 995 120 1005
rect 40 975 50 995
rect 70 985 120 995
rect 145 1090 210 1110
rect 70 975 80 985
rect 40 965 80 975
rect 0 925 40 945
rect 20 755 40 925
rect 145 850 165 1090
rect 185 905 225 915
rect 185 885 195 905
rect 215 885 225 905
rect 185 875 225 885
rect 145 840 185 850
rect 145 820 155 840
rect 175 820 185 840
rect 145 810 185 820
rect 205 755 225 875
rect -50 745 -5 755
rect -50 675 -35 745
rect -15 675 -5 745
rect -50 665 -5 675
rect 20 745 60 755
rect 20 675 30 745
rect 50 675 60 745
rect 20 665 60 675
rect 85 745 125 755
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect 190 745 235 755
rect 190 675 200 745
rect 220 675 235 745
rect 190 665 235 675
rect -50 505 -5 515
rect -50 435 -35 505
rect -15 435 -5 505
rect -50 405 -5 435
rect -50 335 -35 405
rect -15 335 -5 405
rect 40 415 60 665
rect 190 640 210 665
rect 145 620 210 640
rect 145 415 165 620
rect 40 405 100 415
rect 40 395 70 405
rect -50 325 -5 335
rect 60 335 70 395
rect 90 335 100 405
rect 60 325 100 335
rect 125 405 165 415
rect 125 335 135 405
rect 155 335 165 405
rect 125 325 165 335
rect 190 405 235 415
rect 190 335 200 405
rect 220 335 235 405
rect 190 325 235 335
rect 80 290 100 325
rect 80 270 120 290
rect 40 240 80 250
rect 40 230 50 240
rect 0 220 50 230
rect 70 220 80 240
rect 0 210 80 220
rect 0 125 20 210
rect 100 185 120 270
rect 140 255 160 325
rect 140 245 225 255
rect 140 235 195 245
rect 185 225 195 235
rect 215 225 225 245
rect 185 215 225 225
rect 40 175 120 185
rect 40 155 50 175
rect 70 165 120 175
rect 145 175 185 185
rect 70 155 80 165
rect 40 145 80 155
rect 145 155 155 175
rect 175 155 185 175
rect 145 145 185 155
rect 0 105 80 125
rect 60 80 80 105
rect 145 80 165 145
rect -50 70 -5 80
rect -50 0 -35 70
rect -15 0 -5 70
rect -50 -30 -5 0
rect 60 70 100 80
rect 60 0 70 70
rect 90 0 100 70
rect 60 -10 100 0
rect 125 70 165 80
rect 125 0 135 70
rect 155 0 165 70
rect 125 -10 165 0
rect 190 70 235 80
rect 190 0 200 70
rect 220 0 235 70
rect 190 -10 235 0
rect -50 -100 -35 -30
rect -15 -100 -5 -30
rect -50 -110 -5 -100
rect 20 -160 60 -150
rect 20 -230 30 -160
rect 50 -230 60 -160
rect 20 -240 60 -230
rect 125 -160 165 -150
rect 125 -230 135 -160
rect 155 -230 165 -160
rect 125 -240 165 -230
rect -50 -270 235 -260
rect -50 -280 -15 -270
rect -25 -290 -15 -280
rect 5 -280 90 -270
rect 5 -290 15 -280
rect -25 -295 15 -290
rect 80 -290 90 -280
rect 110 -280 235 -270
rect 110 -290 120 -280
rect 80 -295 120 -290
<< viali >>
rect 30 1270 50 1340
rect 135 1270 155 1340
rect 95 1140 115 1210
rect 95 675 115 745
rect -35 435 -15 505
rect -35 335 -15 405
rect 200 335 220 405
rect -35 0 -15 70
rect 200 0 220 70
rect -35 -100 -15 -30
rect 30 -230 50 -160
rect 135 -230 155 -160
<< metal1 >>
rect -50 1340 235 1355
rect -50 1270 30 1340
rect 50 1270 135 1340
rect 155 1270 235 1340
rect -50 1255 235 1270
rect 85 1210 125 1255
rect 85 1140 95 1210
rect 115 1140 125 1210
rect 85 745 125 1140
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect -50 405 -5 435
rect -50 335 -35 405
rect -15 335 -5 405
rect -50 70 -5 335
rect -50 0 -35 70
rect -15 0 -5 70
rect -50 -30 -5 0
rect -50 -100 -35 -30
rect -15 -100 -5 -30
rect -50 -145 -5 -100
rect 190 405 235 415
rect 190 335 200 405
rect 220 335 235 405
rect 190 70 235 335
rect 190 0 200 70
rect 220 0 235 70
rect 190 -145 235 0
rect -50 -160 235 -145
rect -50 -230 30 -160
rect 50 -230 135 -160
rect 155 -230 235 -160
rect -50 -245 235 -230
<< labels >>
rlabel locali 235 710 235 710 3 Q
rlabel locali -50 710 -50 710 7 D
rlabel metal1 -50 -200 -50 -200 7 VN
rlabel locali -50 -270 -50 -270 7 CLK
rlabel locali 235 1175 235 1175 3 Qn
rlabel locali -50 1175 -50 1175 7 Dn
rlabel metal1 -50 1310 -50 1310 7 VP
<< end >>
