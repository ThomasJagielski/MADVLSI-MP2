magic
tech sky130A
timestamp 1614660924
<< nwell >>
rect -70 640 270 1390
<< nmos >>
rect 0 420 15 520
rect 40 420 55 520
rect 105 420 135 520
rect 185 420 200 520
rect 0 -70 15 30
rect 40 -70 55 30
rect 105 -70 135 30
rect 185 -70 200 30
<< pmos >>
rect 0 1140 15 1240
rect 65 1140 80 1240
rect 130 1140 145 1240
rect 185 1140 200 1240
rect 0 660 15 760
rect 65 660 80 760
rect 130 660 145 760
rect 185 660 200 760
<< ndiff >>
rect -50 505 0 520
rect -50 435 -35 505
rect -15 435 0 505
rect -50 420 0 435
rect 15 420 40 520
rect 55 505 105 520
rect 55 435 70 505
rect 90 435 105 505
rect 55 420 105 435
rect 135 505 185 520
rect 135 435 150 505
rect 170 435 185 505
rect 135 420 185 435
rect 200 505 250 520
rect 200 435 215 505
rect 235 435 250 505
rect 200 420 250 435
rect -50 15 0 30
rect -50 -55 -35 15
rect -15 -55 0 15
rect -50 -70 0 -55
rect 15 -70 40 30
rect 55 15 105 30
rect 55 -55 70 15
rect 90 -55 105 15
rect 55 -70 105 -55
rect 135 15 185 30
rect 135 -55 150 15
rect 170 -55 185 15
rect 135 -70 185 -55
rect 200 15 250 30
rect 200 -55 215 15
rect 235 -55 250 15
rect 200 -70 250 -55
<< pdiff >>
rect -50 1225 0 1240
rect -50 1155 -35 1225
rect -15 1155 0 1225
rect -50 1140 0 1155
rect 15 1225 65 1240
rect 15 1155 30 1225
rect 50 1155 65 1225
rect 15 1140 65 1155
rect 80 1225 130 1240
rect 80 1155 95 1225
rect 115 1155 130 1225
rect 80 1140 130 1155
rect 145 1140 185 1240
rect 200 1225 250 1240
rect 200 1155 215 1225
rect 235 1155 250 1225
rect 200 1140 250 1155
rect -50 745 0 760
rect -50 675 -35 745
rect -15 675 0 745
rect -50 660 0 675
rect 15 745 65 760
rect 15 675 30 745
rect 50 675 65 745
rect 15 660 65 675
rect 80 745 130 760
rect 80 675 95 745
rect 115 675 130 745
rect 80 660 130 675
rect 145 660 185 760
rect 200 745 250 760
rect 200 675 215 745
rect 235 675 250 745
rect 200 660 250 675
<< ndiffc >>
rect -35 435 -15 505
rect 70 435 90 505
rect 150 435 170 505
rect 215 435 235 505
rect -35 -55 -15 15
rect 70 -55 90 15
rect 150 -55 170 15
rect 215 -55 235 15
<< pdiffc >>
rect -35 1155 -15 1225
rect 30 1155 50 1225
rect 95 1155 115 1225
rect 215 1155 235 1225
rect -35 675 -15 745
rect 30 675 50 745
rect 95 675 115 745
rect 215 675 235 745
<< psubdiff >>
rect 15 -115 65 -100
rect 15 -185 30 -115
rect 50 -185 65 -115
rect 15 -200 65 -185
rect 135 -115 185 -100
rect 135 -185 150 -115
rect 170 -185 185 -115
rect 135 -200 185 -185
<< nsubdiff >>
rect 15 1355 65 1370
rect 15 1285 30 1355
rect 50 1285 65 1355
rect 15 1270 65 1285
rect 145 1355 195 1370
rect 145 1285 160 1355
rect 180 1285 195 1355
rect 145 1270 195 1285
<< psubdiffcont >>
rect 30 -185 50 -115
rect 150 -185 170 -115
<< nsubdiffcont >>
rect 30 1285 50 1355
rect 160 1285 180 1355
<< poly >>
rect 0 1240 15 1255
rect 65 1240 80 1255
rect 130 1240 145 1255
rect 185 1240 200 1255
rect 0 955 15 1140
rect 65 1085 80 1140
rect 130 1130 145 1140
rect 40 1075 80 1085
rect 40 1055 50 1075
rect 70 1055 80 1075
rect 40 1045 80 1055
rect 105 1115 145 1130
rect 185 1130 200 1140
rect 185 1115 215 1130
rect 40 1010 80 1020
rect 40 990 50 1010
rect 70 990 80 1010
rect 40 980 80 990
rect 0 940 40 955
rect 25 790 40 940
rect 0 775 40 790
rect 0 760 15 775
rect 65 760 80 980
rect 105 785 120 1115
rect 200 915 215 1115
rect 200 905 240 915
rect 200 885 210 905
rect 230 885 240 905
rect 200 875 240 885
rect 160 840 200 850
rect 160 820 170 840
rect 190 820 200 840
rect 160 810 200 820
rect 105 770 145 785
rect 130 760 145 770
rect 185 760 200 810
rect 0 520 15 660
rect 65 650 80 660
rect 130 650 145 660
rect 40 635 80 650
rect 105 635 145 650
rect 40 520 55 635
rect 105 535 120 635
rect 105 520 135 535
rect 185 520 200 660
rect 0 235 15 420
rect 40 365 55 420
rect 40 355 80 365
rect 40 335 50 355
rect 70 335 80 355
rect 40 325 80 335
rect 40 290 80 300
rect 40 270 50 290
rect 70 270 80 290
rect 40 260 80 270
rect 0 220 40 235
rect 25 95 40 220
rect 0 80 40 95
rect 0 30 15 80
rect 65 55 80 260
rect 40 40 80 55
rect 40 30 55 40
rect 105 30 135 420
rect 185 190 200 420
rect 185 180 240 190
rect 185 160 210 180
rect 230 160 240 180
rect 185 150 240 160
rect 160 115 200 125
rect 160 95 170 115
rect 190 95 200 115
rect 160 85 200 95
rect 185 30 200 85
rect 0 -215 15 -70
rect 40 -85 55 -70
rect 105 -215 135 -70
rect 185 -85 200 -70
rect -25 -225 15 -215
rect -25 -245 -15 -225
rect 5 -245 15 -225
rect -25 -255 15 -245
rect 80 -225 135 -215
rect 80 -245 90 -225
rect 110 -245 135 -225
rect 80 -255 135 -245
<< polycont >>
rect 50 1055 70 1075
rect 50 990 70 1010
rect 210 885 230 905
rect 170 820 190 840
rect 50 335 70 355
rect 50 270 70 290
rect 210 160 230 180
rect 170 95 190 115
rect -15 -245 5 -225
rect 90 -245 110 -225
<< locali >>
rect 20 1355 60 1365
rect 20 1285 30 1355
rect 50 1285 60 1355
rect 20 1275 60 1285
rect 150 1355 190 1365
rect 150 1285 160 1355
rect 180 1285 190 1355
rect 150 1275 190 1285
rect -50 1225 -5 1235
rect -50 1155 -35 1225
rect -15 1155 -5 1225
rect -50 1145 -5 1155
rect 20 1225 60 1235
rect 20 1155 30 1225
rect 50 1155 60 1225
rect 20 1145 60 1155
rect 85 1225 125 1235
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 1145 125 1155
rect 205 1225 250 1235
rect 205 1155 215 1225
rect 235 1155 250 1225
rect 205 1145 250 1155
rect 40 1125 60 1145
rect 205 1125 225 1145
rect 40 1105 120 1125
rect 40 1075 80 1085
rect 40 1065 50 1075
rect 0 1055 50 1065
rect 70 1055 80 1075
rect 0 1045 80 1055
rect 0 960 20 1045
rect 100 1020 120 1105
rect 40 1010 120 1020
rect 40 990 50 1010
rect 70 1000 120 1010
rect 160 1105 225 1125
rect 70 990 80 1000
rect 40 980 80 990
rect 0 940 40 960
rect 20 755 40 940
rect 160 850 180 1105
rect 200 905 240 915
rect 200 885 210 905
rect 230 885 240 905
rect 200 875 240 885
rect 160 840 200 850
rect 160 820 170 840
rect 190 820 200 840
rect 160 810 200 820
rect 220 755 240 875
rect -50 745 -5 755
rect -50 675 -35 745
rect -15 675 -5 745
rect -50 665 -5 675
rect 20 745 60 755
rect 20 675 30 745
rect 50 675 60 745
rect 20 665 60 675
rect 85 745 125 755
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect 205 745 250 755
rect 205 675 215 745
rect 235 675 250 745
rect 205 665 250 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect 40 515 60 665
rect 205 635 225 665
rect 160 615 225 635
rect 160 515 180 615
rect 40 505 100 515
rect 40 495 70 505
rect -50 425 -5 435
rect 60 435 70 495
rect 90 435 100 505
rect 60 425 100 435
rect 140 505 180 515
rect 140 435 150 505
rect 170 435 180 505
rect 140 425 180 435
rect 205 505 250 515
rect 205 435 215 505
rect 235 435 250 505
rect 205 425 250 435
rect 80 405 100 425
rect 80 385 120 405
rect 40 355 80 365
rect 40 345 50 355
rect 0 335 50 345
rect 70 335 80 355
rect 0 325 80 335
rect 0 240 20 325
rect 100 300 120 385
rect 40 290 120 300
rect 40 270 50 290
rect 70 280 120 290
rect 70 270 80 280
rect 40 260 80 270
rect 0 220 80 240
rect 60 25 80 220
rect 160 125 180 425
rect 200 180 240 190
rect 200 160 210 180
rect 230 160 240 180
rect 200 150 240 160
rect 160 115 200 125
rect 160 95 170 115
rect 190 95 200 115
rect 160 85 200 95
rect 220 65 240 150
rect 160 45 240 65
rect 160 25 180 45
rect -50 15 -5 25
rect -50 -55 -35 15
rect -15 -55 -5 15
rect -50 -70 -5 -55
rect 60 15 100 25
rect 60 -55 70 15
rect 90 -55 100 15
rect 60 -65 100 -55
rect 140 15 180 25
rect 140 -55 150 15
rect 170 -55 180 15
rect 140 -65 180 -55
rect 205 15 250 25
rect 205 -55 215 15
rect 235 -55 250 15
rect 205 -65 250 -55
rect 20 -115 60 -105
rect 20 -185 30 -115
rect 50 -185 60 -115
rect 20 -195 60 -185
rect 140 -115 180 -105
rect 140 -185 150 -115
rect 170 -185 180 -115
rect 140 -195 180 -185
rect -50 -225 250 -215
rect -50 -235 -15 -225
rect -25 -245 -15 -235
rect 5 -235 90 -225
rect 5 -245 15 -235
rect -25 -255 15 -245
rect 80 -245 90 -235
rect 110 -235 250 -225
rect 110 -245 120 -235
rect 80 -255 120 -245
<< viali >>
rect 30 1285 50 1355
rect 160 1285 180 1355
rect 95 1155 115 1225
rect 95 675 115 745
rect -35 435 -15 505
rect 215 435 235 505
rect -35 -55 -15 15
rect 215 -55 235 15
rect 30 -185 50 -115
rect 150 -185 170 -115
<< metal1 >>
rect -50 1355 250 1370
rect -50 1285 30 1355
rect 50 1285 160 1355
rect 180 1285 250 1355
rect -50 1270 250 1285
rect 85 1225 125 1270
rect 85 1155 95 1225
rect 115 1155 125 1225
rect 85 745 125 1155
rect 85 675 95 745
rect 115 675 125 745
rect 85 665 125 675
rect -50 505 -5 520
rect -50 435 -35 505
rect -15 435 -5 505
rect -50 15 -5 435
rect -50 -55 -35 15
rect -15 -55 -5 15
rect -50 -100 -5 -55
rect 205 505 250 515
rect 205 435 215 505
rect 235 435 250 505
rect 205 15 250 435
rect 205 -55 215 15
rect 235 -55 250 15
rect 205 -100 250 -55
rect -50 -115 250 -100
rect -50 -185 30 -115
rect 50 -185 150 -115
rect 170 -185 250 -115
rect -50 -200 250 -185
<< labels >>
rlabel locali -50 710 -50 710 7 D
port 2 w
rlabel locali -50 1190 -50 1190 7 Dn
port 1 w
rlabel metal1 -50 1325 -50 1325 7 VP
port 6 w
rlabel metal1 -50 -155 -50 -155 7 VN
port 7 w
rlabel locali -50 -225 -50 -225 7 CLK
port 5 w
rlabel locali 250 1190 250 1190 3 Qn
port 3 e
rlabel locali 250 710 250 710 3 Q
port 4 e
<< end >>
