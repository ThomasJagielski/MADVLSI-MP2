magic
tech sky130A
timestamp 1614649743
<< nwell >>
rect -70 705 85 1455
<< nmos >>
rect 0 170 15 270
<< pmos >>
rect 0 1205 15 1305
rect 0 875 15 975
<< ndiff >>
rect -50 255 0 270
rect -50 185 -35 255
rect -15 185 0 255
rect -50 170 0 185
rect 15 255 65 270
rect 15 185 30 255
rect 50 185 65 255
rect 15 170 65 185
<< pdiff >>
rect -50 1290 0 1305
rect -50 1220 -35 1290
rect -15 1220 0 1290
rect -50 1205 0 1220
rect 15 1290 65 1305
rect 15 1220 30 1290
rect 50 1220 65 1290
rect 15 1205 65 1220
rect -50 960 0 975
rect -50 890 -35 960
rect -15 890 0 960
rect -50 875 0 890
rect 15 960 65 975
rect 15 890 30 960
rect 50 890 65 960
rect 15 875 65 890
<< ndiffc >>
rect -35 185 -15 255
rect 30 185 50 255
<< pdiffc >>
rect -35 1220 -15 1290
rect 30 1220 50 1290
rect -35 890 -15 960
rect 30 890 50 960
<< psubdiff >>
rect -50 -50 0 -35
rect -50 -120 -35 -50
rect -15 -120 0 -50
rect -50 -135 0 -120
<< nsubdiff >>
rect -50 1420 0 1435
rect -50 1350 -35 1420
rect -15 1350 0 1420
rect -50 1335 0 1350
<< psubdiffcont >>
rect -35 -120 -15 -50
<< nsubdiffcont >>
rect -35 1350 -15 1420
<< poly >>
rect 0 1305 15 1320
rect 0 1120 15 1205
rect -45 1110 15 1120
rect -45 1090 -35 1110
rect -15 1090 15 1110
rect -45 1080 15 1090
rect 0 975 15 1080
rect 0 865 15 875
rect -45 850 15 865
rect -45 690 -30 850
rect -45 680 35 690
rect -45 675 5 680
rect -45 295 -30 675
rect -5 660 5 675
rect 25 660 35 680
rect -5 650 35 660
rect -45 280 15 295
rect 0 270 15 280
rect 0 155 15 170
<< polycont >>
rect -35 1090 -15 1110
rect 5 660 25 680
<< locali >>
rect -45 1420 -5 1430
rect -45 1350 -35 1420
rect -15 1350 -5 1420
rect -45 1340 -5 1350
rect -45 1290 -5 1300
rect -45 1220 -35 1290
rect -15 1220 -5 1290
rect -45 1210 -5 1220
rect 20 1290 65 1300
rect 20 1220 30 1290
rect 50 1220 65 1290
rect 20 1210 65 1220
rect -50 1110 -5 1120
rect -50 1090 -35 1110
rect -15 1090 -5 1110
rect -50 1080 -5 1090
rect 20 970 40 1210
rect -45 960 -5 970
rect -45 890 -35 960
rect -15 890 -5 960
rect -45 880 -5 890
rect 20 960 60 970
rect 20 890 30 960
rect 50 890 60 960
rect 20 885 60 890
rect 20 860 40 885
rect -45 840 40 860
rect -45 305 -25 840
rect 15 760 65 780
rect 15 690 35 760
rect -5 680 35 690
rect -5 660 5 680
rect 25 660 35 680
rect -5 650 35 660
rect -45 285 40 305
rect 20 265 40 285
rect -45 255 -5 265
rect -45 185 -35 255
rect -15 185 -5 255
rect -45 175 -5 185
rect 20 255 60 265
rect 20 185 30 255
rect 50 185 60 255
rect 20 175 60 185
rect -45 -50 -5 -40
rect -45 -120 -35 -50
rect -15 -120 -5 -50
rect -45 -130 -5 -120
rect -50 -170 65 -150
<< viali >>
rect -35 1350 -15 1420
rect -35 1220 -15 1290
rect -35 890 -15 960
rect -35 185 -15 255
rect -35 -120 -15 -50
<< metal1 >>
rect -50 1420 65 1435
rect -50 1350 -35 1420
rect -15 1350 65 1420
rect -50 1335 65 1350
rect -45 1290 -5 1335
rect -45 1220 -35 1290
rect -15 1220 -5 1290
rect -45 960 -5 1220
rect -45 890 -35 960
rect -15 890 -5 960
rect -45 880 -5 890
rect -45 255 -5 265
rect -45 185 -35 255
rect -15 185 -5 255
rect -45 -35 -5 185
rect -50 -50 65 -35
rect -50 -120 -35 -50
rect -15 -120 65 -50
rect -50 -135 65 -120
<< labels >>
rlabel metal1 -50 1385 -50 1385 7 VP
port 3 w
rlabel locali 65 1255 65 1255 3 Y
port 2 e
rlabel locali 65 770 65 770 3 Ao
port 6 e
rlabel locali -50 1100 -50 1100 7 A
port 1 w
rlabel metal1 -50 -85 -50 -85 7 VN
port 4 w
rlabel locali -50 -160 -50 -160 7 CLK
port 5 w
<< end >>
