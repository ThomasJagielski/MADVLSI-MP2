* SPICE3 file created from D_latch_lvs.ext - technology: sky130A


* Top level circuit D_latch_lvs

X0 a_30_840# CLK VN VN sky130_fd_pr__nfet_01v8 ad=2.5e+11p pd=2.5e+06u as=2e+12p ps=1.2e+07u w=1e+06u l=150000u
X1 VP a_30_1320# a_30_2280# VP sky130_fd_pr__pfet_01v8 ad=1e+12p pd=6e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X2 a_290_1320# CLK VP VP sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=150000u
X3 Q Qn a_290_1320# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_30_1320# CLK D VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X5 a_30_2280# a_30_1320# a_30_n140# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=2.5e+11p ps=2.5e+06u w=1e+06u l=150000u
X6 Qn CLK a_30_2280# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=300000u
X7 Q CLK a_30_1320# VN sky130_fd_pr__nfet_01v8 ad=5e+11p pd=3e+06u as=5e+11p ps=3e+06u w=1e+06u l=300000u
X8 a_290_2280# CLK VP VP sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=150000u
X9 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 VP a_30_2280# a_30_1320# VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_30_n140# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X12 Qn Q a_290_2280# VP sky130_fd_pr__pfet_01v8 ad=5e+11p pd=3e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_30_2280# CLK Dn VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=5e+11p ps=3e+06u w=1e+06u l=150000u
X14 a_30_1320# a_30_2280# a_30_840# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X15 VN Qn Q VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.end

