* SPICE3 file created from CSRL_D_FF.ext - technology: sky130A

X0 a_30_1940# CLK Dn VP sky130_fd_pr__pfet_01v8 ad=2e+08p pd=395000u as=0p ps=0u w=1e+06u l=150000u
X1 Q CLK a_30_1310# VN sky130_fd_pr__nfet_01v8 ad=-2.5e+07p pd=0u as=-4.53743e+16p ps=1.1042e+08u w=1e+06u l=150000u
X2 a_30_0# CLK VN VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=3.35544e+15p ps=0u w=1.9e+06u l=150000u
X3 Qn Q a_290_1940# VP sky130_fd_pr__pfet_01v8 ad=1.20189e+14p pd=0u as=0p ps=0u w=1e+06u l=150000u
X4 VP a_30_1310# a_30_1940# VP sky130_fd_pr__pfet_01v8 ad=-2.5e+07p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 VN Q Qn VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_290_1310# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=150000u
X7 Qn CLK a_30_1940# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_30_1310# CLK D VP sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 VN Qn Q VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=150000u
X10 a_30_1310# a_30_1940# a_30_720# VN sky130_fd_pr__nfet_01v8 ad=-0p pd=0u as=-2.5e+07p ps=1.63445e+08u w=1.9e+06u l=150000u
X11 a_30_1940# a_30_1310# a_30_0# VN sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.9e+06u l=150000u
X12 a_290_1940# CLK VP VP sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=-0p ps=0u w=1e+06u l=150000u
X13 Q Qn a_290_1310# VP sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_30_720# CLK VN VN sky130_fd_pr__nfet_01v8 ad=-0p pd=0u as=0p ps=0u w=1.9e+06u l=150000u
X15 VP a_30_1940# a_30_1310# VP sky130_fd_pr__pfet_01v8 ad=-0p pd=0u as=-0p ps=0u w=1e+06u l=150000u
