magic
tech sky130A
timestamp 1614216702
<< nwell >>
rect -70 635 255 1225
<< nmos >>
rect 0 360 15 550
rect 40 360 55 550
rect 105 450 120 550
rect 170 450 185 550
rect 0 0 15 190
rect 40 0 55 190
rect 105 0 120 100
rect 170 0 185 100
<< pmos >>
rect 0 970 15 1070
rect 65 970 80 1070
rect 130 970 145 1070
rect 170 970 185 1070
rect 0 655 15 755
rect 65 655 80 755
rect 130 655 145 755
rect 170 655 185 755
<< ndiff >>
rect -50 535 0 550
rect -50 465 -35 535
rect -15 465 0 535
rect -50 445 0 465
rect -50 375 -35 445
rect -15 375 0 445
rect -50 360 0 375
rect 15 360 40 550
rect 55 535 105 550
rect 55 465 70 535
rect 90 465 105 535
rect 55 450 105 465
rect 120 535 170 550
rect 120 465 135 535
rect 155 465 170 535
rect 120 450 170 465
rect 185 535 235 550
rect 185 465 200 535
rect 220 465 235 535
rect 185 450 235 465
rect 55 360 80 450
rect -50 175 0 190
rect -50 105 -35 175
rect -15 105 0 175
rect -50 85 0 105
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
rect 15 0 40 190
rect 55 100 80 190
rect 55 85 105 100
rect 55 15 70 85
rect 90 15 105 85
rect 55 0 105 15
rect 120 85 170 100
rect 120 15 135 85
rect 155 15 170 85
rect 120 0 170 15
rect 185 85 235 100
rect 185 15 200 85
rect 220 15 235 85
rect 185 0 235 15
<< pdiff >>
rect -50 1055 0 1070
rect -50 985 -35 1055
rect -15 985 0 1055
rect -50 970 0 985
rect 15 1055 65 1070
rect 15 985 30 1055
rect 50 985 65 1055
rect 15 970 65 985
rect 80 1055 130 1070
rect 80 985 95 1055
rect 115 985 130 1055
rect 80 970 130 985
rect 145 970 170 1070
rect 185 1055 235 1070
rect 185 985 200 1055
rect 220 985 235 1055
rect 185 970 235 985
rect -50 740 0 755
rect -50 670 -35 740
rect -15 670 0 740
rect -50 655 0 670
rect 15 740 65 755
rect 15 670 30 740
rect 50 670 65 740
rect 15 655 65 670
rect 80 740 130 755
rect 80 670 95 740
rect 115 670 130 740
rect 80 655 130 670
rect 145 655 170 755
rect 185 740 235 755
rect 185 670 200 740
rect 220 670 235 740
rect 185 655 235 670
<< ndiffc >>
rect -35 465 -15 535
rect -35 375 -15 445
rect 70 465 90 535
rect 135 465 155 535
rect 200 465 220 535
rect -35 105 -15 175
rect -35 15 -15 85
rect 70 15 90 85
rect 135 15 155 85
rect 200 15 220 85
<< pdiffc >>
rect -35 985 -15 1055
rect 30 985 50 1055
rect 95 985 115 1055
rect 200 985 220 1055
rect -35 670 -15 740
rect 30 670 50 740
rect 95 670 115 740
rect 200 670 220 740
<< psubdiff >>
rect 15 -45 65 -30
rect 15 -115 30 -45
rect 50 -115 65 -45
rect 15 -130 65 -115
rect 120 -45 170 -30
rect 120 -115 135 -45
rect 155 -115 170 -45
rect 120 -130 170 -115
<< nsubdiff >>
rect 15 1185 65 1200
rect 15 1115 30 1185
rect 50 1115 65 1185
rect 15 1100 65 1115
rect 120 1185 170 1200
rect 120 1115 135 1185
rect 155 1115 170 1185
rect 120 1100 170 1115
<< psubdiffcont >>
rect 30 -115 50 -45
rect 135 -115 155 -45
<< nsubdiffcont >>
rect 30 1115 50 1185
rect 135 1115 155 1185
<< poly >>
rect 0 1070 15 1085
rect 65 1070 80 1085
rect 130 1070 145 1085
rect 170 1070 185 1085
rect 0 755 15 970
rect 65 915 80 970
rect 130 960 145 970
rect 40 905 80 915
rect 40 885 50 905
rect 70 885 80 905
rect 40 875 80 885
rect 105 945 145 960
rect 40 840 80 850
rect 40 820 50 840
rect 70 820 80 840
rect 40 810 80 820
rect 65 755 80 810
rect 105 780 120 945
rect 170 915 185 970
rect 145 905 185 915
rect 145 885 155 905
rect 175 885 185 905
rect 145 875 185 885
rect 170 840 225 850
rect 170 820 195 840
rect 215 820 225 840
rect 170 810 225 820
rect 105 765 145 780
rect 130 755 145 765
rect 170 755 185 810
rect 0 550 15 655
rect 65 645 80 655
rect 130 645 145 655
rect 40 630 80 645
rect 105 630 145 645
rect 40 550 55 630
rect 105 550 120 630
rect 170 550 185 655
rect 0 190 15 360
rect 40 350 55 360
rect 40 340 80 350
rect 40 320 50 340
rect 70 320 80 340
rect 40 310 80 320
rect 40 275 80 285
rect 40 255 50 275
rect 70 255 80 275
rect 40 245 80 255
rect 40 190 55 245
rect 105 100 120 450
rect 170 435 185 450
rect 145 420 185 435
rect 145 190 160 420
rect 185 245 225 255
rect 185 225 195 245
rect 215 225 225 245
rect 185 215 225 225
rect 145 180 185 190
rect 145 160 155 180
rect 175 160 185 180
rect 145 150 185 160
rect 210 125 225 215
rect 170 110 225 125
rect 170 100 185 110
rect 0 -145 15 0
rect 40 -15 55 0
rect 105 -145 120 0
rect 170 -15 185 0
rect -25 -155 15 -145
rect -25 -175 -15 -155
rect 5 -175 15 -155
rect -25 -185 15 -175
rect 80 -155 120 -145
rect 80 -175 90 -155
rect 110 -175 120 -155
rect 80 -185 120 -175
<< polycont >>
rect 50 885 70 905
rect 50 820 70 840
rect 155 885 175 905
rect 195 820 215 840
rect 50 320 70 340
rect 50 255 70 275
rect 195 225 215 245
rect 155 160 175 180
rect -15 -175 5 -155
rect 90 -175 110 -155
<< locali >>
rect 20 1185 60 1195
rect 20 1115 30 1185
rect 50 1115 60 1185
rect 20 1105 60 1115
rect 125 1185 165 1195
rect 125 1115 135 1185
rect 155 1115 165 1185
rect 125 1105 165 1115
rect -50 1055 -5 1065
rect -50 985 -35 1055
rect -15 985 -5 1055
rect -50 975 -5 985
rect 20 1055 60 1065
rect 20 985 30 1055
rect 50 985 60 1055
rect 20 975 60 985
rect 85 1055 125 1065
rect 85 985 95 1055
rect 115 985 125 1055
rect 85 975 125 985
rect 190 1055 235 1065
rect 190 985 200 1055
rect 220 985 235 1055
rect 190 975 235 985
rect 40 955 60 975
rect 40 935 120 955
rect 40 905 80 915
rect 40 895 50 905
rect -25 885 50 895
rect 70 885 80 905
rect -25 875 80 885
rect -25 790 -5 875
rect 100 850 120 935
rect 40 840 120 850
rect 40 820 50 840
rect 70 830 120 840
rect 145 905 185 915
rect 145 885 155 905
rect 175 885 185 905
rect 145 875 185 885
rect 70 820 80 830
rect 40 810 80 820
rect -25 770 40 790
rect 20 750 40 770
rect 145 750 165 875
rect 205 850 225 975
rect 185 840 225 850
rect 185 820 195 840
rect 215 820 225 840
rect 185 810 225 820
rect -50 740 -5 750
rect -50 670 -35 740
rect -15 670 -5 740
rect -50 660 -5 670
rect 20 740 60 750
rect 20 670 30 740
rect 50 670 60 740
rect 20 660 60 670
rect 85 740 125 750
rect 85 670 95 740
rect 115 670 125 740
rect 145 740 235 750
rect 145 730 200 740
rect 85 660 125 670
rect 190 670 200 730
rect 220 670 235 740
rect 190 660 235 670
rect 40 545 60 660
rect 190 635 210 660
rect 145 615 210 635
rect 145 545 165 615
rect -50 535 -5 545
rect -50 465 -35 535
rect -15 465 -5 535
rect 40 535 100 545
rect 40 525 70 535
rect -50 445 -5 465
rect 60 465 70 525
rect 90 465 100 535
rect 60 455 100 465
rect 125 535 165 545
rect 125 465 135 535
rect 155 465 165 535
rect 125 455 165 465
rect 190 535 235 545
rect 190 465 200 535
rect 220 465 235 535
rect 190 455 235 465
rect -50 375 -35 445
rect -15 375 -5 445
rect -50 365 -5 375
rect 80 390 100 455
rect 80 370 120 390
rect 40 340 80 350
rect 40 330 50 340
rect 0 320 50 330
rect 70 320 80 340
rect 0 310 80 320
rect 0 225 20 310
rect 100 285 120 370
rect 40 275 120 285
rect 40 255 50 275
rect 70 265 120 275
rect 70 255 80 265
rect 40 245 80 255
rect 140 255 160 455
rect 140 245 225 255
rect 140 235 195 245
rect 185 225 195 235
rect 215 225 225 245
rect 0 205 35 225
rect 185 215 225 225
rect -50 175 -5 185
rect -50 105 -35 175
rect -15 105 -5 175
rect -50 85 -5 105
rect -50 15 -35 85
rect -15 15 -5 85
rect 15 95 35 205
rect 145 180 185 190
rect 145 160 155 180
rect 175 160 185 180
rect 145 150 185 160
rect 145 95 165 150
rect 15 85 100 95
rect 15 75 70 85
rect -50 5 -5 15
rect 60 15 70 75
rect 90 15 100 85
rect 60 5 100 15
rect 125 85 165 95
rect 125 15 135 85
rect 155 15 165 85
rect 125 5 165 15
rect 190 85 235 95
rect 190 15 200 85
rect 220 15 235 85
rect 190 5 235 15
rect 20 -45 60 -35
rect 20 -115 30 -45
rect 50 -115 60 -45
rect 20 -125 60 -115
rect 125 -45 165 -35
rect 125 -115 135 -45
rect 155 -115 165 -45
rect 125 -125 165 -115
rect -50 -155 235 -145
rect -50 -165 -15 -155
rect -25 -175 -15 -165
rect 5 -165 90 -155
rect 5 -175 15 -165
rect -25 -185 15 -175
rect 80 -175 90 -165
rect 110 -165 235 -155
rect 110 -175 120 -165
rect 80 -185 120 -175
<< viali >>
rect 30 1115 50 1185
rect 135 1115 155 1185
rect 95 985 115 1055
rect 95 670 115 740
rect -35 465 -15 535
rect 200 465 220 535
rect -35 375 -15 445
rect -35 105 -15 175
rect -35 15 -15 85
rect 200 15 220 85
rect 30 -115 50 -45
rect 135 -115 155 -45
<< metal1 >>
rect -50 1185 235 1200
rect -50 1115 30 1185
rect 50 1115 135 1185
rect 155 1115 235 1185
rect -50 1100 235 1115
rect 85 1055 125 1100
rect 85 985 95 1055
rect 115 985 125 1055
rect 85 740 125 985
rect 85 670 95 740
rect 115 670 125 740
rect 85 660 125 670
rect -50 535 -5 545
rect -50 465 -35 535
rect -15 465 -5 535
rect -50 445 -5 465
rect -50 375 -35 445
rect -15 375 -5 445
rect -50 175 -5 375
rect -50 105 -35 175
rect -15 105 -5 175
rect -50 85 -5 105
rect -50 15 -35 85
rect -15 15 -5 85
rect -50 -30 -5 15
rect 190 535 235 545
rect 190 465 200 535
rect 220 465 235 535
rect 190 85 235 465
rect 190 15 200 85
rect 220 15 235 85
rect 190 -30 235 15
rect -50 -45 235 -30
rect -50 -115 30 -45
rect 50 -115 135 -45
rect 155 -115 235 -45
rect -50 -130 235 -115
<< labels >>
rlabel metal1 -50 -85 -50 -85 7 VN
rlabel locali -50 -155 -50 -155 7 CLK
rlabel metal1 -50 1155 -50 1155 7 VP
rlabel locali -50 1020 -50 1020 7 Dn
rlabel locali -50 705 -50 705 7 D
rlabel locali 235 705 235 705 3 Q
rlabel locali 235 1020 235 1020 3 Qn
<< end >>
